/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 958;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_322d746c,
        64'h75616665_642d6972,
        64'h742c786e_6c780074,
        64'h6c756166_65642d69,
        64'h72742c78_6e6c7800,
        64'h6c617564_2d73692c,
        64'h786e6c78_00746e65,
        64'h73657270_2d747075,
        64'h72726574_6e692c78,
        64'h6e6c7800_68746469,
        64'h772d326f_6970672c,
        64'h786e6c78_00687464,
        64'h69772d6f_6970672c,
        64'h786e6c78_00322d74,
        64'h6c756166_65642d74,
        64'h756f642c_786e6c78,
        64'h00746c75_61666564,
        64'h2d74756f_642c786e,
        64'h6c780032_2d737475,
        64'h706e692d_6c6c612c,
        64'h786e6c78_00737475,
        64'h706e692d_6c6c612c,
        64'h786e6c78_0072656c,
        64'h6c6f7274_6e6f632d,
        64'h6f697067_00736c6c,
        64'h65632d6f_69706723,
        64'h00737365_72646461,
        64'h2d63616d_2d6c6163,
        64'h6f6c0070_772d656c,
        64'h62617369_64007365,
        64'h676e6172_2d656761,
        64'h746c6f76_0079636e,
        64'h65757165_72662d78,
        64'h616d2d69_7073006f,
        64'h69746172_2d6b6373,
        64'h2c786e6c_78007374,
        64'h69622d72_6566736e,
        64'h6172742d_6d756e2c,
        64'h786e6c78_00737469,
        64'h622d7373_2d6d756e,
        64'h2c786e6c_78007473,
        64'h6978652d_6f666966,
        64'h2c786e6c_7800796c,
        64'h696d6166_2c786e6c,
        64'h7800736b_636f6c63,
        64'h0073656d_616e2d6b,
        64'h636f6c63_00656461,
        64'h72672d64_65657073,
        64'h00687464_69772d6f,
        64'h692d6765_72007466,
        64'h6968732d_67657200,
        64'h73747075_72726574,
        64'h6e690074_6e657261,
        64'h702d7470_75727265,
        64'h746e6900_64656570,
        64'h732d746e_65727275,
        64'h63007665_646e2c76,
        64'h63736972_00797469,
        64'h726f6972_702d7861,
        64'h6d2c7663_73697200,
        64'h73656d61_6e2d6765,
        64'h72006465_646e6574,
        64'h78652d73_74707572,
        64'h7265746e_69007365,
        64'h676e6172_0073656d,
        64'h616e2d74_75707475,
        64'h6f2d6b63_6f6c6300,
        64'h736c6c65_632d6b63,
        64'h6f6c6323_00646564,
        64'h6e657073_75732d65,
        64'h74617473_2d6e6961,
        64'h74657200_72656767,
        64'h6972742d_746c7561,
        64'h6665642c_78756e69,
        64'h6c00736f_69706700,
        64'h656c646e_61687000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_00736c6c,
        64'h65632d74_70757272,
        64'h65746e69_23007469,
        64'h6c70732d_626c7400,
        64'h65707974_2d756d6d,
        64'h00617369_2c766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745f65_63697665,
        64'h64007963_6e657571,
        64'h6572662d_6b636f6c,
        64'h63007963_6e657571,
        64'h6572662d_65736162,
        64'h656d6974_00687461,
        64'h702d7475_6f647473,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'hb5000000_04000000,
        64'h03000000_ffffffff,
        64'hfe020000_04000000,
        64'h03000000_ffffffff,
        64'hed020000_04000000,
        64'h03000000_01000000,
        64'he0020000_04000000,
        64'h03000000_00000000,
        64'hc9020000_04000000,
        64'h03000000_08000000,
        64'hb8020000_04000000,
        64'h03000000_08000000,
        64'ha8020000_04000000,
        64'h03000000_00000000,
        64'h94020000_04000000,
        64'h03000000_00000000,
        64'h82020000_04000000,
        64'h03000000_00000000,
        64'h70020000_04000000,
        64'h03000000_00000000,
        64'h60020000_04000000,
        64'h03000000_00000100,
        64'h00000000_00000040,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h50020000_00000000,
        64'h03000000_00000000,
        64'h612e3030_2e312d6f,
        64'h6970672d_7370782c,
        64'h786e6c78_1b000000,
        64'h15000000_03000000,
        64'h02000000_44020000,
        64'h04000000_03000000,
        64'h00000030_30303030,
        64'h30303440_6f697067,
        64'h01000000_02000000,
        64'h00800000_00000000,
        64'h00000030_00000000,
        64'h67000000_10000000,
        64'h03000000_00007fe3,
        64'h023e1800_32020000,
        64'h06000000_03000000,
        64'h00000000_03000000,
        64'h72010000_08000000,
        64'h03000000_03000000,
        64'h61010000_04000000,
        64'h03000000_006b726f,
        64'h7774656e_5b000000,
        64'h08000000_03000000,
        64'h00687465_2d637369,
        64'h72776f6c_1b000000,
        64'h0c000000_03000000,
        64'h00000000_30303030,
        64'h30303033_40687465,
        64'h2d637369_72776f6c,
        64'h01000000_02000000,
        64'h02000000_27020000,
        64'h00000000_03000000,
        64'he40c0000_e40c0000,
        64'h18020000_08000000,
        64'h03000000_20bcbe00,
        64'h06020000_04000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00000000,
        64'h746f6c73_2d697073,
        64'h2d636d6d_1b000000,
        64'h0d000000_03000000,
        64'h00000030_40636d6d,
        64'h01000000_04000000,
        64'hf7010000_04000000,
        64'h03000000_08000000,
        64'he0010000_04000000,
        64'h03000000_01000000,
        64'hcf010000_04000000,
        64'h03000000_01000000,
        64'hbf010000_04000000,
        64'h03000000_00377865,
        64'h746e696b_b3010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000020_00000000,
        64'h67000000_10000000,
        64'h03000000_02000000,
        64'h02000000_72010000,
        64'h08000000_03000000,
        64'h03000000_61010000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00612e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_00622e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h1b000000_28000000,
        64'h03000000_00000000,
        64'h30303030_30303032,
        64'h40697073_2d737078,
        64'h01000000_02000000,
        64'h00100000_00000000,
        64'h00000019_00000000,
        64'h67000000_10000000,
        64'h03000000_00000062,
        64'h66726570_61702c72,
        64'h65706170_1b000000,
        64'h0e000000_03000000,
        64'h00003030_30303030,
        64'h39314072_65706170,
        64'h01000000_02000000,
        64'h006c6f72_746e6f63,
        64'h2b010000_08000000,
        64'h03000000_03000000,
        64'h61010000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000018,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h07000000_06000000,
        64'h05000000_04000000,
        64'h72010000_10000000,
        64'h03000000_00007265,
        64'h6d69745f_6270612c,
        64'h706c7570_1b000000,
        64'h0f000000_03000000,
        64'h00003030_30303030,
        64'h38314072_656d6974,
        64'h01000000_02000000,
        64'h00003774_756f5f6b,
        64'h6c630036_74756f5f,
        64'h6b6c6300_3574756f,
        64'h5f6b6c63_00347475,
        64'h6f5f6b6c_63003374,
        64'h756f5f6b_6c630032,
        64'h74756f5f_6b6c6300,
        64'h3174756f_5f6b6c63,
        64'hfd000000_3f000000,
        64'h03000000_00000000,
        64'h05000000_00000000,
        64'h04000000_ac010000,
        64'h10000000_03000000,
        64'h00006b6c_63615f69,
        64'h78615f73_00316e69,
        64'h5f6b6c63_a0010000,
        64'h13000000_03000000,
        64'h01000000_94010000,
        64'h04000000_03000000,
        64'h00000000_6472617a,
        64'h69772d67_6e696b63,
        64'h6f6c632c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_00100000,
        64'h00000000_00000017,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h01000000_f0000000,
        64'h04000000_03000000,
        64'h00000000_30303030,
        64'h30303731_40726f74,
        64'h6172656e_65672d6b,
        64'h636f6c63_01000000,
        64'h02000000_04000000,
        64'h87010000_04000000,
        64'h03000000_02000000,
        64'h7d010000_04000000,
        64'h03000000_01000000,
        64'h72010000_04000000,
        64'h03000000_03000000,
        64'h61010000_04000000,
        64'h03000000_00c20100,
        64'h53010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_2b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_17010000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_48010000,
        64'h04000000_03000000,
        64'h07000000_35010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_17010000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_2b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_17010000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'h10010000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'h05000000_b5000000,
        64'h04000000_03000000,
        64'h006b6c63_5f697861,
        64'hfd000000_08000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_01000000,
        64'hf0000000_04000000,
        64'h03000000_006b636f,
        64'h6c632d64_65786966,
        64'h1b000000_0c000000,
        64'h03000000_006b6c63,
        64'h5f697861_01000000,
        64'h02000000_04000000,
        64'hb5000000_04000000,
        64'h03000000_006b6c63,
        64'h5f666572_fd000000,
        64'h08000000_03000000,
        64'h00c2eb0b_4b000000,
        64'h04000000_03000000,
        64'h01000000_f0000000,
        64'h04000000_03000000,
        64'h006b636f_6c632d64,
        64'h65786966_1b000000,
        64'h0c000000_03000000,
        64'h006b6c63_5f666572,
        64'h01000000_0000736b,
        64'h636f6c63_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha40b0000_11030000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'hdc0b0000_38000000,
        64'hed0e0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_a0018402,
        64'h13058593_00000597,
        64'h01f41413_0010041b,
        64'he911d05f_f0ef057e,
        64'h65a14505_ebcff0ef,
        64'h04050513_00001517,
        64'he84ff0ef_e4060805,
        64'h05132005_85931141,
        64'h02faf537_65f1b38d,
        64'hee0ff0ef_35450513,
        64'h00001517_bbd90ae5,
        64'h05130000_1517f78f,
        64'hf0ef8526_efcff0ef,
        64'h1b050513_00001517,
        64'hf08ff0ef_1a450513,
        64'h00001517_bbfd0d65,
        64'h05130000_1517fa0f,
        64'hf0ef8526_f24ff0ef,
        64'h1d850513_00001517,
        64'hf30ff0ef_1cc50513,
        64'h00001517_c92984aa,
        64'hc3dff0ef_8556865e,
        64'h020b2583_f4cff0ef,
        64'h3a850513_00001517,
        64'hf3849de3_08090913,
        64'h080a0993_f64ff0ef,
        64'h248512a5_05130000,
        64'h1517ff3a_1be383bf,
        64'hf0ef0a05_000a4503,
        64'hf80ff0ef_3cc50513,
        64'h00001517_80fff0ef,
        64'h01093503_f94ff0ef,
        64'h3d050513_00001517,
        64'h823ff0ef_00893503,
        64'hfa8ff0ef_3d450513,
        64'h00001517_837ff0ef,
        64'hfb898a13_00093503,
        64'hfc0ff0ef_3dc50513,
        64'h00001517_ff2a1be3,
        64'h895ff0ef_0a05000a,
        64'h4503f909_8a13fdef,
        64'hf0ef3da5_05130000,
        64'h1517ff9a_19e38b3f,
        64'hf0ef0a05_0007c503,
        64'h014d07b3_4a01ffef,
        64'hf0eff809_8d133de5,
        64'h05130000_15178d3f,
        64'hf0ef0ff4_f513817f,
        64'hf0ef3da5_05130000,
        64'h15174c11_4cc11005,
        64'h1b630201_09130801,
        64'h099384aa_8b0ad33f,
        64'hf0ef850a_46057101,
        64'h04892583_845ff0ef,
        64'h20850513_00001517,
        64'h893ff0ef_4556857f,
        64'hf0ef3fa5_05130000,
        64'h15178a5f_f0ef4546,
        64'h869ff0ef_3ec50513,
        64'h00001517_8f7ff0ef,
        64'h652687bf_f0ef3de5,
        64'h05130000_1517909f,
        64'hf0ef7502_88dff0ef,
        64'h3e050513_00001517,
        64'h91bff0ef_656289ff,
        64'hf0ef3da5_05130000,
        64'h15178edf_f0ef4552,
        64'h8b1ff0ef_3dc50513,
        64'h00001517_8ffff0ef,
        64'h45428c3f_f0ef3de5,
        64'h05130000_1517911f,
        64'hf0ef4532_8d5ff0ef,
        64'h3e050513_00001517,
        64'h923ff0ef_45228e7f,
        64'hf0ef3e25_05130000,
        64'h1517975f_f0ef6502,
        64'h8f9ff0ef_3e450513,
        64'h00001517_905ff0ef,
        64'h3d050513_00001517,
        64'hbf5154f9_915ff0ef,
        64'h2d850513_00001517,
        64'h9a3ff0ef_8526927f,
        64'hf0ef3da5_05130000,
        64'h1517933f_f0ef3ce5,
        64'h05130000_1517c905,
        64'h84aa890a_e41ff0ef,
        64'h850a4585_46057101,
        64'h951ff0ef_3d450513,
        64'h00001517_80826125,
        64'h6d026ca2_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_64468526,
        64'h60e6fa04_011354fd,
        64'h981ff0ef_3dc50513,
        64'h00001517_c90ddeff,
        64'hf0ef8bae_8aaa1080,
        64'he06ae466_e862f05a,
        64'hf852fc4e_e0cae4a6,
        64'hec86ec5e_f456e8a2,
        64'h711db765_54798082,
        64'h61696baa_6b4a6aea,
        64'h7a0a79aa_794a74ea,
        64'h640e60ae_8522547d,
        64'h9d1ff0ef_40450513,
        64'h00001517_c5dff0ef,
        64'hc61ff0ef_c65ff0ef,
        64'hc69ff0ef_c6dff0ef,
        64'hc71ff0ef_c75ff0ef,
        64'hc79ff0ef_a805c7ff,
        64'hf0efc8bf_f0ef4531,
        64'h45814605_4401f930,
        64'h46e32004_849319fd,
        64'ha19ff0ef_46c50513,
        64'h00001517_e7990369,
        64'he7b30689_1c639041,
        64'h29011442_8c49cb7f,
        64'hf0ef9041_03051413,
        64'h0085151b_cc5ff0ef,
        64'hfc941ae3_04040413,
        64'hff7a17e3_892af15f,
        64'hf0ef0a05_854a0007,
        64'hc5830144_07b30400,
        64'h0b934a01_c69ff0ef,
        64'h850a0400_05938622,
        64'h4901ff55_1ee3cfff,
        64'hf0efe004_84133e80,
        64'h0b130fe0_0a93e951,
        64'h20048493_d1dff0ef,
        64'h454985a2_0ff67613,
        64'h00166613_0015161b,
        64'hf4dff0ef_0ff47593,
        64'hf55ff0ef_0ff5f593,
        64'h0084559b_f61ff0ef,
        64'h0ff5f593_0104559b,
        64'hf6dff0ef_45010184,
        64'h559bfee7_9be30785,
        64'h00c68023_00f106b3,
        64'h08000713_567d4781,
        64'h0209d993_842e84aa,
        64'he55ee95a_ed56f152,
        64'hf94ae586_fd26e1a2,
        64'h02061993_f54e7155,
        64'h80829141_15428d3d,
        64'h8ff90057_979b1701,
        64'h67090107_d79b0105,
        64'h179b4105_551b0105,
        64'h151b8d2d_00c59513,
        64'h8da9893d_0045d51b,
        64'h8da99141_15428d5d,
        64'h05220085_579b8082,
        64'h07f57513_8d2d0045,
        64'h15938d2d_8d3d0045,
        64'hd51b0075_d79b8de9,
        64'h80820141_853e6402,
        64'h60a257f5_e1114781,
        64'hf89ff0ef_c51157f9,
        64'hefbff0ef_c91157fd,
        64'heb7ff0ef_fc6de07f,
        64'hf0ef347d_4429b8ff,
        64'hf0ef5aa5_05130000,
        64'h1517c89f_f0efe022,
        64'he4061141_80826105,
        64'h00153513_64a26442,
        64'h60e20004_051bfc94,
        64'h0ce3e3bf_f0efeb3f,
        64'hf0ef5d25_05130000,
        64'h151785aa_842ae57f,
        64'hf0ef0290_05134000,
        64'h05b70770_0613fbdf,
        64'hf0ef4485_e822ec06,
        64'he4261101_80820141,
        64'h00153513_157d6402,
        64'h60a20004_051bef3f,
        64'hf0ef60c5_051385a2,
        64'h00001517_e8dff0ef,
        64'h842ae9bf_f0efe022,
        64'he4060370_05134581,
        64'h06500613_11418082,
        64'h61056902_64a26442,
        64'h60e20015_3513f565,
        64'h05130004_051b0124,
        64'h986388bd_00f91b63,
        64'h45014785_ecdff0ef,
        64'hed1ff0ef_842aed7f,
        64'hf0ef84aa_eddff0ef,
        64'hee1ff0ef_ee5ff0ef,
        64'h892aef3f_f0efe04a,
        64'he426e822_ec064521,
        64'h1aa00593_08700613,
        64'h1101bfcd_45018082,
        64'h61056902_64a26442,
        64'h60e24505_f89ff0ef,
        64'h458569a5_05130000,
        64'h1517fe99_15e3c00d,
        64'hf29ff0ef_892a347d,
        64'hf39ff0ef_45014581,
        64'h09500613_44857104,
        64'h0413e04a_ec06e426,
        64'h6409e822_1101ccff,
        64'hf06f6105_69450513,
        64'h00001517_60e26442,
        64'hda5ff0ef_852e65a2,
        64'hce9ff0ef_6dc50513,
        64'h00001517_cf5ff0ef,
        64'h8522cfbf_f0efe42e,
        64'hec066e25_05130000,
        64'h1517842a_e8221101,
        64'h80826145_64e27402,
        64'h70a2f47d_147d0007,
        64'hd4634187_d79b0185,
        64'h179bfabf_f0efeb5f,
        64'hf0ef8532_06400413,
        64'h6622ec1f_f0ef0ff4,
        64'h7513ec9f_f0ef0ff5,
        64'h75130084_551bed5f,
        64'hf0ef0ff5_75130104,
        64'h551bee1f_f0ef0184,
        64'h551bee9f_f0ef0404,
        64'he513febf_f0ef84aa,
        64'h842eec26_f022e432,
        64'hf4067179_f03ff06f,
        64'h0ff00513_8082557d,
        64'hb7d900d7_00230785,
        64'h00f60733_06c82683,
        64'hff698b05_5178b77d,
        64'hd6b80785_00074703,
        64'h00f50733_80824501,
        64'hd3b84719_dbb8577d,
        64'h200007b7_02b6e163,
        64'h0007869b_20000837,
        64'h20000537_fff58b85,
        64'h537c2000_0737d3b8,
        64'h200007b7_10600713,
        64'hfff537fd_00010320,
        64'h079304b7_61630007,
        64'h871b4781_200006b7,
        64'hdbb85779_200007b7,
        64'h06b7ee63_10000793,
        64'h80826105_64a2d3b8,
        64'h4719dbb8_644260e2,
        64'h0ff47513_577d2000,
        64'h07b7e23f_f0ef7e65,
        64'h05130000_1517eb1f,
        64'hf0ef9101_15024088,
        64'he39ff0ef_80450513,
        64'h00002517_e3958b85,
        64'h240153fc_57e0ff65,
        64'h8b050647_849353f8,
        64'hd3b81060_07132000,
        64'h07b7fff5_37fd0001,
        64'h06400793_d7a8dbb8,
        64'h5779e426_e822ec06,
        64'h200007b7_1101e7ff,
        64'hf06f6105_83450513,
        64'h00002517_64a260e2,
        64'h6442d03c_4799e97f,
        64'hf0ef85a5_05130000,
        64'h2517f25f_f0ef9101,
        64'h02049513_2481eaff,
        64'hf0ef8525_05130000,
        64'h25175064_d03c1660,
        64'h0793ec3f_f0ef8865,
        64'h05130000_2517f51f,
        64'hf0ef9101_02049513,
        64'h2481edbf_f0ef87e5,
        64'h05130000_25175064,
        64'hd03c1040_07932000,
        64'h0437fff5_37fd0001,
        64'h47a9c3b8_47292000,
        64'h07b7f03f_f0efe426,
        64'he822ec06_89e50513,
        64'h11010000_25178082,
        64'h25014108_8082c10c,
        64'h80826105_60e2ecff,
        64'hf0ef0091_4503ed7f,
        64'hf0ef0081_4503f55f,
        64'hf0efec06_002c1101,
        64'h80826145_694264e2,
        64'h740270a2_fe9410e3,
        64'hef9ff0ef_00914503,
        64'hf01ff0ef_34610081,
        64'h4503f81f_f0ef0ff5,
        64'h7513002c_00895533,
        64'h54e10380_0413892a,
        64'hf406e84a_ec26f022,
        64'h71798082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f3bf_f0ef0091,
        64'h4503f43f_f0ef3461,
        64'h00814503_fc3ff0ef,
        64'h0ff57513_002c0089,
        64'h553b54e1_4461892a,
        64'hf406e84a_ec26f022,
        64'h71798082_00f58023,
        64'h0007c783_00e580a3,
        64'h97aa8111_00074703,
        64'h973e00f5_771396e7,
        64'h87930000_1797b7f5,
        64'h0405f93f_f0ef8082,
        64'h01416402_60a2e509,
        64'h00044503_842ae406,
        64'he0221141_808200e7,
        64'h88230200_071300e7,
        64'h8423fc70_071300e7,
        64'h8623470d_00a78223,
        64'h0ff57513_00e78023,
        64'h0085551b_0ff57713,
        64'h00e78623_f8000713,
        64'h00078223_100007b7,
        64'h02b5553b_0045959b,
        64'h808200a7_0023dfe5,
        64'h0207f793_01474783,
        64'h10000737_80820205,
        64'h75130147_c5031000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_b8458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h27f000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
